<svg aria-hidden="true" style="position:absolute;width:0;height:0;overflow:hidden" xmlns="http://www.w3.org/2000/svg">
  <defs>
    <symbol id="icon-close-iscon" viewBox="0 0 32 32">
<path d="M32 3.721l-3.721-3.721-12.279 12.279-12.279-12.279-3.721 3.721 12.279 12.279-12.279 12.279 3.721 3.721 12.279-12.279 12.279 12.279 3.721-3.721-12.279-12.279 12.279-12.279z"></path>
</symbol>
<symbol id="icon-menu-icon" viewBox="0 0 32 32">
<path stroke-linejoin="round" stroke-linecap="round" stroke-miterlimit="4" stroke-width="3.3333" d="M2 20.667h28M2 11.333h28"></path>
</symbol>
<symbol id="icon-facebook-icon" viewBox="0 0 32 32">
<path d="M32 16.040c0-8.854-7.168-16.040-16-16.040s-16 7.186-16 16.040c0 7.763 5.504 14.228 12.8 15.719v-10.907h-3.2v-4.812h3.2v-4.010c0-3.096 2.512-5.614 5.6-5.614h4v4.812h-3.2c-0.88 0-1.6 0.722-1.6 1.604v3.208h4.8v4.812h-4.8v11.148c8.080-0.802 14.4-7.635 14.4-15.96z"></path>
</symbol>
<symbol id="icon-youtube-icon" viewBox="0 0 32 32">
<path d="M18.672 15.722l-3.743-1.747c-0.327-0.152-0.595 0.018-0.595 0.38v3.29c0 0.362 0.268 0.532 0.595 0.38l3.742-1.747c0.328-0.153 0.328-0.403 0.002-0.557zM16 0c-8.837 0-16 7.163-16 16s7.163 16 16 16c8.837 0 16-7.163 16-16s-7.163-16-16-16zM16 22.5c-8.19 0-8.333-0.738-8.333-6.5s0.143-6.5 8.333-6.5c8.19 0 8.333 0.738 8.333 6.5s-0.143 6.5-8.333 6.5z"></path>
</symbol>
<symbol id="icon-instagram-icon" viewBox="0 0 32 32">
<path d="M23.385 0h-14.769c-2.284 0.002-4.474 0.911-6.089 2.526s-2.524 3.805-2.526 6.089v14.769c0.002 2.284 0.911 4.474 2.526 6.089s3.805 2.524 6.089 2.526h14.769c2.284-0.003 4.474-0.911 6.089-2.526s2.524-3.805 2.526-6.089v-14.769c-0.003-2.284-0.911-4.474-2.526-6.089s-3.805-2.524-6.089-2.526zM16 23.385c-1.461 0-2.888-0.433-4.103-1.244s-2.161-1.965-2.72-3.314c-0.559-1.349-0.705-2.834-0.42-4.267s0.988-2.748 2.021-3.781c1.033-1.033 2.349-1.736 3.781-2.021s2.917-0.139 4.267 0.42c1.349 0.559 2.503 1.505 3.314 2.72s1.244 2.642 1.244 4.103c-0.002 1.958-0.781 3.835-2.165 5.22s-3.262 2.163-5.22 2.165zM25.231 8.615c-0.365 0-0.722-0.108-1.026-0.311s-0.54-0.491-0.68-0.829c-0.14-0.337-0.176-0.709-0.105-1.067s0.247-0.687 0.505-0.945c0.258-0.258 0.587-0.434 0.945-0.505s0.729-0.035 1.067 0.105c0.337 0.14 0.626 0.376 0.829 0.68s0.311 0.661 0.311 1.026c0 0.49-0.195 0.959-0.541 1.305s-0.816 0.541-1.305 0.541zM20.923 16c0 0.974-0.289 1.926-0.83 2.735s-1.31 1.441-2.209 1.813c-0.9 0.373-1.889 0.47-2.844 0.28s-1.832-0.659-2.521-1.347c-0.688-0.689-1.157-1.566-1.347-2.521s-0.092-1.945 0.28-2.844 1.004-1.668 1.813-2.209c0.81-0.541 1.761-0.83 2.735-0.83 1.306 0 2.558 0.519 3.481 1.442s1.442 2.175 1.442 3.481z"></path>
</symbol>
  </defs>
</svg>